`timescale 1ns/1ps
module snapshot_tb;

  reg clk, rst_n;
  reg left, right, shoot;
  reg enemy_spawn;
  reg [4:0] enemy_init_x;
  reg [3:0] enemy_init_y;

  wire [4:0] player_x;
  wire [3:0] player_y;
  wire [4:0] bullet_x;
  wire [3:0] bullet_y;
  wire        bullet_active;

  wire [4:0] enemy0_x, enemy1_x, enemy2_x;
  wire [3:0] enemy0_y, enemy1_y, enemy2_y;
  wire        enemy0_active, enemy1_active, enemy2_active;

  wire        hit;
  wire [7:0]  hit_count;
  wire [7:0]  score;

  game_design dut(
    .clk(clk), .rst_n(rst_n),
    .left(left), .right(right), .shoot(shoot),
    .enemy_spawn(enemy_spawn), .enemy_init_x(enemy_init_x), .enemy_init_y(enemy_init_y),
    .player_x(player_x), .player_y(player_y),
    .bullet_x(bullet_x), .bullet_y(bullet_y), .bullet_active(bullet_active),
    .enemy0_x(enemy0_x), .enemy0_y(enemy0_y), .enemy0_active(enemy0_active),
    .enemy1_x(enemy1_x), .enemy1_y(enemy1_y), .enemy1_active(enemy1_active),
    .enemy2_x(enemy2_x), .enemy2_y(enemy2_y), .enemy2_active(enemy2_active),
    .hit(hit), .hit_count(hit_count), .score(score)
  );

  initial begin clk = 0; forever #1 clk = ~clk; end

  integer cycle;
  initial begin
    $dumpfile("snapshot.vcd");
    $dumpvars(0, snapshot_tb);

    left=0; right=0; shoot=0;
    enemy_spawn=0; enemy_init_x=0; enemy_init_y=0;
    rst_n=0; #5; rst_n=1; #2;
    cycle = 0;

    #(45*2);
    left = 1; #2; left = 0;
    #(9*2);
    shoot = 1; #2; shoot = 0;
    #(12*2);
    left = 1; #2; left = 0;
    #(7*2);
    shoot = 1; #2; shoot = 0;
    #(24*2);
    shoot = 1; #2; shoot = 0;
    #(13*2);
    right = 1; #2; right = 0;
    #(10*2);
    right = 1; #2; right = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(18*2);
    left = 1; #2; left = 0;
    #(9*2);
    right = 1; #2; right = 0;
    #(9*2);
    shoot = 1; #2; shoot = 0;
    #(7*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(27*2);
    shoot = 1; #2; shoot = 0;
    #(7*2);
    left = 1; #2; left = 0;
    #(19*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(10*2);
    right = 1; #2; right = 0;
    #(11*2);
    shoot = 1; #2; shoot = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(38*2);
    shoot = 1; #2; shoot = 0;
    #(6*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(15*2);
    left = 1; #2; left = 0;
    #(12*2);
    shoot = 1; #2; shoot = 0;
    #(31*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(4*2);
    right = 1; #2; right = 0;
    #(8*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(4*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(4*2);
    right = 1; #2; right = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(11*2);
    shoot = 1; #2; shoot = 0;
    #(13*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(10*2);
    shoot = 1; #2; shoot = 0;
    #(20*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(18*2);
    left = 1; #2; left = 0;
    #(7*2);
    shoot = 1; #2; shoot = 0;
    #(19*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(10*2);
    shoot = 1; #2; shoot = 0;
    #(7*2);
    right = 1; #2; right = 0;
    #(4*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(7*2);
    shoot = 1; #2; shoot = 0;
    #(19*2);
    left = 1; #2; left = 0;
    #(6*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(12*2);
    shoot = 1; #2; shoot = 0;
    #(10*2);
    left = 1; #2; left = 0;
    #(7*2);
    left = 1; #2; left = 0;
    #(12*2);
    right = 1; #2; right = 0;
    #(22*2);
    shoot = 1; #2; shoot = 0;
    #(6*2);
    left = 1; #2; left = 0;
    #(18*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(3*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(8*2);
    shoot = 1; #2; shoot = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(4*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(30*2);
    right = 1; #2; right = 0;
    #(7*2);
    right = 1; #2; right = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(19*2);
    left = 1; #2; left = 0;
    #(14*2);
    shoot = 1; #2; shoot = 0;
    #(7*2);
    right = 1; #2; right = 0;
    #(73*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(6*2);
    right = 1; #2; right = 0;
    #(8*2);
    right = 1; #2; right = 0;
    #(13*2);
    right = 1; #2; right = 0;
    #(12*2);
    right = 1; #2; right = 0;
    #(10*2);
    shoot = 1; #2; shoot = 0;
    #(21*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(6*2);
    left = 1; #2; left = 0;
    #(12*2);
    left = 1; #2; left = 0;
    #(5*2);
    shoot = 1; #2; shoot = 0;
    #(10*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(4*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(5*2);
    left = 1; #2; left = 0;
    #(7*2);
    shoot = 1; #2; shoot = 0;
    #(14*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(4*2);
    right = 1; #2; right = 0;
    #(9*2);
    right = 1; #2; right = 0;
    #(5*2);
    right = 1; #2; right = 0;
    #(2000*2);
    $finish;
  end
endmodule
